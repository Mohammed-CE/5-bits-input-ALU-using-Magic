magic
tech scmos
timestamp 1607580023
<< error_p >>
rect 776 3576 778 3580
<< error_s >>
rect -248 6312 -246 6313
rect 1274 6308 1275 6314
rect 2030 6309 2031 6315
<< metal1 >>
rect -1117 6392 -1113 6396
rect -537 6392 -533 6396
rect 223 6392 227 6396
rect 983 6392 987 6396
rect 1739 6392 1743 6396
rect 2495 6392 2499 6396
rect -1281 6184 -1277 6188
rect -1281 5860 -1277 5864
rect -1281 5536 -1277 5540
rect -1281 5216 -1277 5220
rect -1281 4900 -1277 4904
rect -1300 -92 -1296 4420
rect -1292 -80 -1288 4432
rect -1284 -68 -1280 4444
rect -1276 -56 -1272 4456
rect -1268 -44 -1264 4468
rect -1021 4424 -1017 4577
rect -297 4436 -293 4565
rect 451 4448 455 4576
rect 1255 4460 1259 4564
rect 2207 4472 2211 4552
rect -1048 -8 -1044 3880
rect -1040 1796 -1036 3868
rect -100 3796 -96 3880
rect -992 3728 -988 3732
rect -992 3532 -988 3536
rect -616 3404 -612 3408
rect -1040 436 -1036 1792
rect -1032 1328 -1028 3396
rect -1032 340 -1028 1324
rect -1024 1288 -1020 3356
rect -964 3220 -960 3224
rect -964 3024 -960 3028
rect -1024 244 -1020 1284
rect -1016 820 -1012 2888
rect -1016 148 -1012 816
rect -1008 780 -1004 2848
rect -1008 52 -1004 776
rect -1000 596 -996 2664
rect -1000 484 -996 592
rect -992 692 -988 2760
rect -968 2712 -964 2716
rect 120 2457 124 2628
rect 132 2465 136 3108
rect 144 2473 148 3136
rect 156 2481 160 3616
rect 168 2489 172 3644
rect 508 3576 775 3580
rect 508 3466 512 3576
rect 516 3474 520 3568
rect 524 3482 528 3560
rect 532 3490 536 3552
rect 540 3498 544 3532
rect 540 3494 547 3498
rect 532 3486 547 3490
rect 524 3478 547 3482
rect 647 3474 656 3478
rect 516 3470 547 3474
rect 508 3462 547 3466
rect 652 3092 656 3474
rect 500 3088 656 3092
rect 500 2815 504 3088
rect 424 2811 459 2815
rect 500 2811 507 2815
rect 424 2720 428 2811
rect 424 2716 624 2720
rect 168 2485 175 2489
rect 156 2477 173 2481
rect 144 2469 173 2473
rect 132 2461 173 2465
rect 120 2453 173 2457
rect 356 2109 360 2676
rect 392 2316 396 2465
rect 392 2224 396 2312
rect 577 2152 581 2156
rect 477 1892 481 1896
rect 365 1884 369 1888
rect 81 1672 85 1676
rect -411 1288 -407 1292
rect -411 812 -407 816
rect -992 388 -988 688
rect 348 633 358 637
rect 406 568 410 633
rect 620 536 624 2716
rect 660 576 664 3544
rect 680 1112 684 3552
rect 700 1648 704 3560
rect 708 2184 712 3568
rect 776 2720 780 3580
rect 316 532 624 536
rect 180 288 184 308
rect 8 -260 12 -96
rect 20 -252 24 -84
rect 32 -244 36 -72
rect 44 -236 48 -60
rect 56 -228 60 -48
rect 56 -232 61 -228
rect 44 -240 61 -236
rect 32 -248 61 -244
rect 316 -248 320 532
rect 344 520 516 524
rect 344 248 348 520
rect 400 456 406 460
rect 410 456 568 460
rect 368 52 372 268
rect 376 148 380 276
rect 384 176 388 284
rect 392 132 396 292
rect 392 52 396 128
rect 400 68 404 300
rect 392 48 400 52
rect 508 24 512 48
rect 564 24 568 456
rect 744 436 748 2608
rect 752 340 756 2064
rect 760 288 764 1532
rect 768 280 772 992
rect 776 784 780 2628
rect 776 700 780 780
rect 784 1912 788 2444
rect 784 1376 788 1908
rect 784 840 788 1372
rect 776 272 780 460
rect 784 304 788 836
rect 792 2016 796 2548
rect 792 1480 796 2012
rect 792 944 796 1476
rect 792 408 796 940
rect 792 388 796 404
rect 804 1920 808 2452
rect 804 1384 808 1916
rect 804 848 808 1380
rect 852 1324 856 3108
rect 860 1856 864 3136
rect 868 2388 872 3616
rect 876 2924 880 3644
rect 2536 3548 2540 4784
rect 2544 3556 2548 5100
rect 2552 3564 2556 5420
rect 2564 3572 2568 5744
rect 2572 3580 2576 6068
rect 2536 3020 2540 3060
rect 2544 3048 2548 3060
rect 876 2820 880 2920
rect 1016 2772 1020 2776
rect 868 2296 872 2384
rect 924 2336 928 2500
rect 1016 2236 1020 2240
rect 860 1752 864 1852
rect 924 1800 928 1964
rect 1016 1700 1020 1704
rect 852 1224 856 1320
rect 924 1264 928 1428
rect 1016 1164 1020 1168
rect 804 312 808 844
rect 924 728 928 892
rect 1016 628 1020 632
rect 924 296 928 356
rect 508 -8 512 20
rect 760 -44 764 128
rect 768 -56 772 56
rect 800 4 804 192
rect 752 -252 756 -96
rect 776 -132 780 -84
rect 800 -188 804 0
rect 808 -92 812 96
rect 20 -256 61 -252
rect 8 -264 61 -260
rect 808 -284 812 -96
rect 816 68 820 144
rect 824 136 828 144
rect 816 64 824 68
rect 816 -52 820 64
rect 816 -56 824 -52
rect 816 -124 820 -56
rect 816 -128 824 -124
rect 816 -244 820 -128
rect 816 -248 824 -244
<< metal2 >>
rect -956 6384 -952 6388
rect -246 6310 -242 6316
rect 514 6309 518 6315
rect 1274 6308 1278 6314
rect 2030 6309 2034 6315
rect 2286 6304 2290 6310
rect 2786 6308 2790 6314
rect -1000 6097 -990 6101
rect 2363 6072 2576 6076
rect 2363 5748 2568 5752
rect 2363 5424 2556 5428
rect 2363 5104 2548 5108
rect 2523 4856 2540 4860
rect 2363 4788 2540 4792
rect -1264 4468 2207 4472
rect -1272 4456 1255 4460
rect 1259 4456 1264 4460
rect -1280 4444 451 4448
rect 455 4444 462 4448
rect -1288 4432 -297 4436
rect -293 4432 -288 4436
rect -1296 4420 -1021 4424
rect -1017 4420 -1013 4424
rect -1044 3880 -100 3884
rect -1036 3868 -616 3872
rect -1087 3728 -996 3732
rect -400 3644 168 3648
rect 172 3644 876 3648
rect -400 3616 156 3620
rect 160 3616 868 3620
rect 784 3576 2572 3580
rect 520 3568 708 3572
rect 712 3568 2564 3572
rect 528 3560 700 3564
rect 704 3560 2552 3564
rect 536 3552 680 3556
rect 684 3552 2544 3556
rect 664 3544 2536 3548
rect -1087 3532 -996 3536
rect 544 3532 660 3536
rect 547 3522 551 3526
rect 547 3426 551 3430
rect -1028 3396 -616 3400
rect -1020 3356 -588 3360
rect -1087 3220 -968 3224
rect -372 3136 144 3140
rect 148 3136 860 3140
rect -372 3108 132 3112
rect 136 3108 852 3112
rect 957 3052 3036 3056
rect -1087 3024 -968 3028
rect 880 2920 896 2924
rect -1012 2888 -588 2892
rect 599 2859 603 2863
rect -1004 2848 -592 2852
rect 880 2816 896 2820
rect -60 2808 -56 2812
rect 599 2811 648 2815
rect -988 2760 -944 2764
rect 599 2763 603 2767
rect -1087 2712 -972 2716
rect 644 2676 648 2811
rect 780 2716 896 2720
rect 364 2672 648 2676
rect -996 2664 -944 2668
rect -376 2628 120 2632
rect 124 2628 776 2632
rect 748 2608 896 2612
rect 736 2548 792 2552
rect 796 2548 816 2552
rect -976 2532 -968 2536
rect 736 2517 740 2548
rect 267 2513 740 2517
rect 273 2465 392 2469
rect 760 2452 804 2456
rect 808 2452 816 2456
rect 760 2421 764 2452
rect 788 2444 812 2448
rect 269 2417 764 2421
rect 872 2384 896 2388
rect 396 2312 453 2316
rect 872 2292 896 2296
rect 396 2220 453 2224
rect 712 2180 896 2184
rect 360 2105 453 2109
rect 756 2064 896 2068
rect 796 2012 816 2016
rect 356 1997 453 2001
rect 356 1824 360 1997
rect 412 1933 416 1937
rect 808 1916 816 1920
rect 788 1908 812 1912
rect 864 1852 896 1856
rect 404 1845 408 1849
rect 356 1820 516 1824
rect -1036 1792 -464 1796
rect -460 1792 -439 1796
rect -1087 1656 -828 1660
rect -824 1656 -816 1660
rect -1087 1460 -828 1464
rect -824 1460 -816 1464
rect -1028 1324 -448 1328
rect -444 1324 -439 1328
rect -1025 1284 -1024 1288
rect -1020 1284 -420 1288
rect -1087 1148 -796 1152
rect -792 1148 -788 1152
rect 469 1148 473 1152
rect -1087 952 -796 956
rect -792 952 -788 956
rect -1012 816 -416 820
rect -1004 776 -424 780
rect -420 776 -415 780
rect 180 740 184 744
rect -988 688 -767 692
rect -1087 640 -800 644
rect -796 640 -792 644
rect 344 637 348 736
rect 498 681 502 685
rect 498 633 502 637
rect -996 592 -767 596
rect 498 585 502 589
rect -996 480 -20 484
rect 28 480 32 484
rect 406 460 410 564
rect 512 528 516 1820
rect 864 1748 896 1752
rect 704 1644 896 1648
rect 764 1532 896 1536
rect 796 1476 816 1480
rect 808 1380 816 1384
rect 788 1372 812 1376
rect 856 1320 896 1324
rect 856 1220 896 1224
rect 684 1108 896 1112
rect 772 992 896 996
rect 796 940 816 944
rect 808 844 816 848
rect 788 836 812 840
rect 780 780 896 784
rect 780 696 896 700
rect 664 572 896 576
rect 780 460 896 464
rect -1036 432 0 436
rect 104 432 744 436
rect 796 404 816 408
rect -988 384 -12 388
rect 24 384 28 388
rect 32 384 792 388
rect -1028 336 0 340
rect 104 336 752 340
rect 184 308 804 312
rect 808 308 817 312
rect 404 300 784 304
rect 788 300 812 304
rect 396 292 924 296
rect 388 284 760 288
rect 380 276 768 280
rect 372 268 776 272
rect -1020 240 0 244
rect 192 240 348 244
rect 188 192 404 196
rect 508 192 800 196
rect 804 192 828 196
rect 104 172 384 176
rect -1012 144 0 148
rect 104 144 376 148
rect 512 144 816 148
rect 820 144 824 148
rect 900 144 904 148
rect 396 128 432 132
rect 764 128 824 132
rect 32 96 404 100
rect 508 96 808 100
rect 812 96 828 100
rect 404 64 432 68
rect 772 56 824 60
rect -1004 48 0 52
rect 104 48 368 52
rect 900 48 904 52
rect 512 20 564 24
rect 32 0 404 4
rect 508 0 800 4
rect 804 0 828 4
rect -1044 -12 508 -8
rect -1264 -48 56 -44
rect 60 -48 760 -44
rect 900 -48 904 -44
rect -1272 -60 44 -56
rect 48 -60 768 -56
rect 780 -64 824 -60
rect 780 -68 784 -64
rect -1280 -72 32 -68
rect 36 -72 784 -68
rect -1288 -84 20 -80
rect 24 -84 776 -80
rect -1296 -96 8 -92
rect 12 -96 752 -92
rect 812 -96 828 -92
rect 780 -136 824 -132
rect 900 -144 904 -140
rect 804 -192 828 -188
rect 68 -200 72 -196
rect 900 -240 904 -236
rect 161 -252 316 -248
rect 756 -256 820 -252
rect 812 -288 828 -284
rect 76 -304 80 -300
<< m2contact >>
rect 2359 6072 2363 6076
rect 2572 6068 2576 6072
rect 2359 5748 2363 5752
rect 2564 5744 2568 5748
rect 2359 5424 2363 5428
rect 2552 5420 2556 5424
rect 2359 5104 2363 5108
rect 2544 5100 2548 5104
rect 2359 4788 2363 4792
rect 2536 4784 2540 4788
rect -1268 4468 -1264 4472
rect -1276 4456 -1272 4460
rect -1284 4444 -1280 4448
rect -1292 4432 -1288 4436
rect -1300 4420 -1296 4424
rect 2207 4468 2211 4472
rect 1255 4456 1259 4460
rect 451 4444 455 4448
rect -297 4432 -293 4436
rect -1021 4420 -1017 4424
rect -1048 3880 -1044 3884
rect -100 3880 -96 3884
rect -1040 3868 -1036 3872
rect -616 3868 -612 3872
rect -996 3728 -992 3732
rect -404 3644 -400 3648
rect 168 3644 172 3648
rect -404 3616 -400 3620
rect 156 3616 160 3620
rect -996 3532 -992 3536
rect -1040 1792 -1036 1796
rect -1040 432 -1036 436
rect -1032 3396 -1028 3400
rect -616 3396 -612 3400
rect -1032 1324 -1028 1328
rect -1032 336 -1028 340
rect -1024 3356 -1020 3360
rect -588 3356 -584 3360
rect -968 3220 -964 3224
rect -376 3136 -372 3140
rect 144 3136 148 3140
rect -376 3108 -372 3112
rect 132 3108 136 3112
rect -968 3024 -964 3028
rect -1024 1284 -1020 1288
rect -1024 240 -1020 244
rect -1016 2888 -1012 2892
rect -588 2888 -584 2892
rect -1016 816 -1012 820
rect -1016 144 -1012 148
rect -1008 2848 -1004 2852
rect -592 2848 -588 2852
rect -992 2760 -988 2764
rect -1008 776 -1004 780
rect -1000 2664 -996 2668
rect -1000 592 -996 596
rect -1000 480 -996 484
rect -972 2712 -968 2716
rect -380 2628 -376 2632
rect 120 2628 124 2632
rect 876 3644 880 3648
rect 868 3616 872 3620
rect 516 3568 520 3572
rect 708 3568 712 3572
rect 524 3560 528 3564
rect 700 3560 704 3564
rect 532 3552 536 3556
rect 680 3552 684 3556
rect 660 3544 664 3548
rect 540 3532 544 3536
rect 360 2672 364 2676
rect 392 2465 396 2469
rect 392 2312 396 2316
rect 453 2312 457 2316
rect 392 2220 396 2224
rect 453 2220 457 2224
rect 356 2105 360 2109
rect 453 2105 457 2109
rect 453 1997 457 2001
rect -439 1792 -435 1796
rect -816 1656 -812 1660
rect -816 1460 -812 1464
rect -439 1324 -435 1328
rect -788 1148 -784 1152
rect -788 952 -784 956
rect -415 776 -411 780
rect -992 688 -988 692
rect -792 640 -788 644
rect 344 633 348 637
rect 406 564 410 568
rect 780 3576 784 3580
rect 860 3136 864 3140
rect 776 2716 780 2720
rect 852 3108 856 3112
rect 776 2628 780 2632
rect 708 2180 712 2184
rect 744 2608 748 2612
rect 700 1644 704 1648
rect 680 1108 684 1112
rect 660 572 664 576
rect 0 432 4 436
rect -992 384 -988 388
rect 0 336 4 340
rect 180 308 184 312
rect 0 240 4 244
rect 0 144 4 148
rect -1008 48 -1004 52
rect 0 48 4 52
rect -1048 -12 -1044 -8
rect -1268 -48 -1264 -44
rect 56 -48 60 -44
rect -1276 -60 -1272 -56
rect 44 -60 48 -56
rect -1284 -72 -1280 -68
rect 32 -72 36 -68
rect -1292 -84 -1288 -80
rect 20 -84 24 -80
rect -1300 -96 -1296 -92
rect 8 -96 12 -92
rect 512 524 516 528
rect 406 456 410 460
rect 400 300 404 304
rect 392 292 396 296
rect 384 284 388 288
rect 376 276 380 280
rect 344 244 348 248
rect 368 268 372 272
rect 384 172 388 176
rect 376 144 380 148
rect 368 48 372 52
rect 392 128 396 132
rect 432 128 436 132
rect 400 64 404 68
rect 432 64 436 68
rect 508 48 512 52
rect 508 20 512 24
rect 744 432 748 436
rect 752 2064 756 2068
rect 752 336 756 340
rect 760 1532 764 1536
rect 760 284 764 288
rect 768 992 772 996
rect 792 2548 796 2552
rect 776 780 780 784
rect 776 696 780 700
rect 784 2444 788 2448
rect 784 1908 788 1912
rect 784 1372 788 1376
rect 784 836 788 840
rect 768 276 772 280
rect 776 460 780 464
rect 792 2012 796 2016
rect 792 1476 796 1480
rect 792 940 796 944
rect 792 404 796 408
rect 792 384 796 388
rect 804 2452 808 2456
rect 804 1916 808 1920
rect 804 1380 808 1384
rect 2572 3576 2576 3580
rect 2564 3568 2568 3572
rect 2552 3560 2556 3564
rect 2544 3552 2548 3556
rect 2536 3544 2540 3548
rect 876 2920 880 2924
rect 896 2920 900 2924
rect 876 2816 880 2820
rect 896 2816 900 2820
rect 896 2716 900 2720
rect 896 2608 900 2612
rect 868 2384 872 2388
rect 896 2384 900 2388
rect 868 2292 872 2296
rect 896 2292 900 2296
rect 896 2180 900 2184
rect 896 2064 900 2068
rect 860 1852 864 1856
rect 896 1852 900 1856
rect 860 1748 864 1752
rect 896 1748 900 1752
rect 896 1644 900 1648
rect 896 1532 900 1536
rect 852 1320 856 1324
rect 896 1320 900 1324
rect 852 1220 856 1224
rect 896 1220 900 1224
rect 896 1108 900 1112
rect 896 992 900 996
rect 804 844 808 848
rect 896 780 900 784
rect 896 696 900 700
rect 896 572 900 576
rect 896 460 900 464
rect 804 308 808 312
rect 784 300 788 304
rect 924 292 928 296
rect 776 268 780 272
rect 800 192 804 196
rect 564 20 568 24
rect 760 128 764 132
rect 508 -12 512 -8
rect 760 -48 764 -44
rect 768 56 772 60
rect 768 -60 772 -56
rect 816 144 820 148
rect 800 0 804 4
rect 776 -84 780 -80
rect 316 -252 320 -248
rect 752 -96 756 -92
rect 776 -136 780 -132
rect 800 -192 804 -188
rect 808 96 812 100
rect 808 -96 812 -92
rect 752 -256 756 -252
rect 824 144 828 148
rect 824 128 828 132
rect 824 56 828 60
rect 824 -64 828 -60
rect 824 -136 828 -132
rect 820 -256 824 -252
rect 808 -288 812 -284
use sm  sm_0
timestamp 1607580023
transform 1 0 824 0 1 96
box 0 -384 80 100
use comparator  comparator_0
timestamp 1607580023
transform 1 0 -815 0 1 556
box 0 0 1284 1248
use sd  sd_0
timestamp 1607580023
transform 1 0 432 0 1 96
box -32 -96 80 100
use notnor  notnor_0
timestamp 1607580023
transform 1 0 0 0 -1 484
box -20 0 192 484
use and2  and2_1
timestamp 1607580023
transform 1 0 462 0 1 609
box -104 -24 36 84
use transmission4  transmission4_1
timestamp 1607580023
transform 1 0 892 0 1 1260
box -80 -424 128 108
use transmission4  transmission4_0
timestamp 1607580023
transform 1 0 892 0 1 724
box -80 -424 128 108
use transmission4  transmission4_2
timestamp 1607580023
transform 1 0 892 0 1 1796
box -80 -424 128 108
use nor  nor_2
timestamp 1605567036
transform 1 0 109 0 1 -240
box -48 -60 52 40
use adder5bit  adder5bit_0
timestamp 1607580023
transform 1 0 -1420 0 1 3508
box 428 -880 1376 368
use and2  and2_0
timestamp 1607580023
transform 1 0 563 0 1 2787
box -104 -24 36 84
use transmission4  transmission4_5
timestamp 1607580023
transform 1 0 449 0 1 2257
box -80 -424 128 108
use transmission4  transmission4_3
timestamp 1607580023
transform 1 0 892 0 1 2332
box -80 -424 128 108
use transmission4  transmission4_4
timestamp 1607580023
transform 1 0 892 0 1 2868
box -80 -424 128 108
use nor  nor_1
timestamp 1605567036
transform 1 0 595 0 1 3486
box -48 -60 52 40
use nor  nor_0
timestamp 1605567036
transform 1 0 221 0 1 2477
box -48 -60 52 40
use multiplayer  multiplayer_0
timestamp 1607580023
transform 1 0 -1273 0 1 6092
box -96 -1584 3800 300
<< labels >>
rlabel metal1 1016 2772 1020 2776 7 o0
rlabel metal1 1016 2236 1020 2240 7 o1
rlabel metal1 1016 1700 1020 1704 7 o2
rlabel metal1 1016 1164 1020 1168 7 o3
rlabel metal1 1016 628 1020 632 7 o4
rlabel metal2 900 144 904 148 1 o5
rlabel metal2 900 48 904 52 1 o6
rlabel metal2 900 -48 904 -44 1 o7
rlabel metal2 900 -144 904 -140 1 o8
rlabel metal2 900 -240 904 -236 1 o9
rlabel metal2 -60 2808 -56 2812 1 cout
rlabel metal1 -964 3220 -960 3224 1 b2
rlabel metal1 -992 3532 -988 3536 1 b1
rlabel metal1 -992 3728 -988 3732 1 b0
rlabel metal2 24 384 28 388 1 vdd
rlabel metal2 28 480 32 484 1 gnd
rlabel m2contact 0 48 4 52 1 a4
rlabel m2contact 0 144 4 148 1 a3
rlabel m2contact 0 240 4 244 1 a2
rlabel m2contact 0 336 4 340 1 a1
rlabel m2contact 0 432 4 436 1 a0
rlabel metal1 392 48 396 52 1 s1
rlabel metal1 400 144 404 148 1 s0
rlabel metal1 -964 3024 -960 3028 1 b3
rlabel metal1 -968 2712 -964 2716 1 b4
rlabel metal2 471 1150 471 1150 1 a<=b
rlabel metal2 180 740 184 744 1 a>=b
rlabel metal2 -458 1794 -458 1794 1 a0
rlabel metal2 -822 1658 -822 1658 1 b0
rlabel metal2 -822 1462 -822 1462 1 b1
rlabel metal2 -442 1326 -442 1326 1 a1
rlabel metal1 -409 1290 -409 1290 1 a2
rlabel metal2 -790 1150 -790 1150 1 b2
rlabel metal2 -790 954 -790 954 1 b3
rlabel metal1 -409 814 -409 814 1 a3
rlabel metal2 -418 778 -418 778 1 a4
rlabel metal2 -794 642 -794 642 1 b4
rlabel metal1 83 1674 83 1674 1 cin
rlabel metal1 2497 6394 2497 6394 5 a0
rlabel metal1 1741 6394 1741 6394 5 a1
rlabel metal1 985 6394 985 6394 5 a2
rlabel metal1 225 6394 225 6394 5 a3
rlabel metal1 -535 6394 -535 6394 5 a4
rlabel metal1 -1279 4902 -1279 4902 1 b4
rlabel metal1 -1280 5218 -1280 5218 1 b3
rlabel metal1 -1280 5538 -1280 5538 1 b2
rlabel metal1 -1280 5862 -1280 5862 1 b1
rlabel metal1 -1280 6186 -1280 6186 1 b0
rlabel metal2 -954 6386 -954 6386 1 gnd
rlabel metal1 -1115 6394 -1115 6394 5 vdd
rlabel metal2 549 3524 549 3524 1 vdd
rlabel metal2 549 3428 549 3428 1 gnd
rlabel metal2 70 -198 70 -198 1 vdd
rlabel metal2 78 -302 78 -302 1 gnd
rlabel metal2 601 2765 601 2765 1 gnd
rlabel metal2 601 2861 601 2861 1 vdd
rlabel metal1 479 1894 479 1894 1 s1
rlabel metal1 367 1886 367 1886 1 s0
rlabel metal1 579 2154 579 2154 1 OZ
rlabel metal2 500 587 500 587 1 gnd
rlabel metal2 500 635 500 635 1 ONEg
rlabel metal2 500 683 500 683 1 vdd
rlabel metal2 414 1935 414 1935 1 vdd
rlabel metal2 406 1847 406 1847 1 gnd
<< end >>
