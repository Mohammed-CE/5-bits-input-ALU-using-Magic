magic
tech scmos
timestamp 1606847121
<< metal1 >>
rect 1072 608 1076 988
rect 1080 612 1084 1016
rect 1072 604 1080 608
rect 1052 596 1080 600
rect 1052 512 1056 596
rect 1180 592 1216 596
rect 1072 588 1080 592
rect 1072 484 1076 588
rect 1080 4 1084 584
rect 1236 568 1252 572
rect 1248 184 1252 568
rect 1092 180 1096 184
<< metal2 >>
rect 592 1016 1080 1020
rect 592 988 1072 992
rect 872 640 1084 644
rect 1176 640 1204 644
rect 904 544 1116 548
rect 1176 544 1204 548
rect 620 508 1052 512
rect 620 480 1072 484
rect 908 228 1100 232
rect 932 180 1088 184
rect 1132 180 1248 184
rect 868 132 1100 136
rect 616 0 1080 4
<< polycontact >>
rect 1216 592 1220 596
rect 1232 568 1236 572
<< m2contact >>
rect 588 1016 592 1020
rect 1080 1016 1084 1020
rect 588 988 592 992
rect 1072 988 1076 992
rect 1176 592 1180 596
rect 616 508 620 512
rect 1052 508 1056 512
rect 616 480 620 484
rect 1072 480 1076 484
rect 1088 180 1092 184
rect 1248 180 1252 184
rect 612 0 616 4
rect 1080 0 1084 4
use adder5bit  adder5bit_0
timestamp 1606847121
transform 1 0 -428 0 1 880
box 428 -880 1376 368
use nor  nor_0
timestamp 1605567036
transform 1 0 1128 0 1 604
box -48 -60 52 40
use or  or_0
timestamp 1606069941
transform 1 0 1204 0 1 544
box 0 0 80 100
use not  not_0
timestamp 1605560378
transform 1 0 1092 0 -1 180
box 4 -52 40 48
<< end >>
