magic
tech scmos
timestamp 1607341315
<< metal1 >>
rect 156 292 160 300
rect 736 292 740 300
rect 1496 292 1500 300
rect 2256 292 2260 300
rect 3012 292 3016 300
rect 3768 292 3772 300
rect -4 92 4 96
rect 156 -32 160 8
rect 340 -28 344 12
rect 736 -32 740 8
rect 748 -32 752 8
rect 996 -32 1000 -16
rect 1496 -32 1500 8
rect 1508 -32 1512 8
rect 1756 -32 1760 -16
rect 2256 -32 2260 8
rect 2268 -32 2272 8
rect 2512 -32 2516 -16
rect 3012 -32 3016 8
rect 3024 -32 3028 8
rect 3628 -20 3632 -12
rect 3268 -32 3272 -20
rect 3768 -32 3772 4
rect 3780 -32 3784 4
rect 340 -36 344 -32
rect -4 -232 4 -228
rect 156 -356 160 -308
rect 340 -352 344 -312
rect 736 -356 740 -316
rect 748 -356 752 -316
rect 996 -356 1000 -340
rect 340 -360 344 -356
rect 1496 -357 1500 -317
rect 1508 -356 1512 -316
rect 1756 -356 1760 -340
rect 2256 -356 2260 -316
rect 2268 -356 2272 -316
rect 2512 -356 2516 -340
rect 3012 -356 3016 -316
rect 3024 -356 3028 -316
rect 3268 -356 3272 -340
rect 3628 -344 3632 -336
rect 3768 -356 3772 -320
rect 3780 -356 3784 -320
rect -4 -556 4 -552
rect 156 -680 160 -632
rect 340 -672 344 -632
rect 340 -680 344 -676
rect 736 -680 740 -640
rect 748 -680 752 -640
rect 996 -676 1000 -664
rect 1496 -676 1500 -635
rect 1508 -676 1512 -636
rect 1756 -676 1760 -664
rect 2256 -676 2260 -636
rect 2268 -676 2272 -636
rect 2512 -676 2516 -664
rect 3012 -676 3016 -636
rect 3024 -676 3028 -636
rect 3268 -676 3272 -664
rect 3628 -668 3632 -660
rect 3768 -676 3772 -640
rect 3780 -676 3784 -640
rect -4 -876 4 -872
rect 156 -992 160 -952
rect 340 -988 344 -956
rect 340 -996 344 -992
rect 736 -996 740 -956
rect 748 -996 752 -956
rect 996 -992 1000 -984
rect 1496 -992 1500 -952
rect 1508 -992 1512 -952
rect 1756 -992 1760 -984
rect 2256 -996 2260 -956
rect 2268 -996 2272 -956
rect 2512 -992 2516 -984
rect 3012 -996 3016 -956
rect 3024 -992 3028 -952
rect 3268 -992 3272 -984
rect 3628 -988 3632 -980
rect 3768 -992 3772 -956
rect 3780 -992 3784 -956
rect -4 -1192 4 -1188
rect 40 -1315 44 -1280
rect 224 -1384 228 -1248
rect 364 -1288 368 -1224
rect 2228 -1260 2232 -1257
rect -80 -1480 -76 -1432
rect 252 -1516 256 -1512
rect 552 -1528 556 -1420
rect 596 -1444 600 -1294
rect 764 -1327 768 -1288
rect 916 -1396 920 -1270
rect 1100 -1300 1104 -1275
rect 1508 -1284 1512 -1267
rect 2228 -1272 2232 -1264
rect 596 -1448 639 -1444
rect 976 -1528 980 -1524
rect 1276 -1580 1280 -1428
rect 1300 -1528 1304 -1352
rect 1356 -1432 1360 -1290
rect 1528 -1340 1532 -1276
rect 1676 -1384 1680 -1274
rect 1860 -1288 1864 -1272
rect 1356 -1436 1380 -1432
rect 1724 -1516 1728 -1512
rect 2016 -1580 2020 -1340
rect 2024 -1540 2028 -1420
rect 2116 -1444 2120 -1285
rect 2236 -1317 2240 -1292
rect 2316 -1328 2320 -1276
rect 2432 -1288 2436 -1275
rect 2684 -1300 2688 -1224
rect 3012 -1277 3016 -1274
rect 2872 -1300 2876 -1283
rect 3052 -1288 3056 -1284
rect 2828 -1428 2832 -1418
rect 2116 -1448 2188 -1444
rect 2828 -1520 2832 -1432
rect 2528 -1528 2532 -1524
rect 2852 -1540 2856 -1352
rect 3024 -1456 3028 -1292
rect 3188 -1343 3192 -1267
rect 3628 -1304 3632 -1296
rect 3268 -1336 3272 -1304
rect 3648 -1312 3652 -1224
rect 3024 -1460 3140 -1456
rect 3796 -1520 3800 -1364
rect 3480 -1540 3484 -1536
<< metal2 >>
rect 240 288 340 292
rect 344 288 748 292
rect 752 288 996 292
rect 1000 288 1508 292
rect 1512 288 1756 292
rect 1760 288 2268 292
rect 2272 288 2512 292
rect 2516 288 3024 292
rect 3028 288 3268 292
rect 3272 288 3780 292
rect 600 -16 996 -12
rect 1360 -16 1756 -12
rect 2120 -16 2512 -12
rect 2876 -20 3268 -16
rect 240 -32 340 -28
rect 600 -340 996 -336
rect 1360 -340 1756 -336
rect 2120 -340 2512 -336
rect 2516 -340 2520 -336
rect 2876 -340 3268 -336
rect 3272 -340 3276 -336
rect 240 -356 340 -352
rect 600 -664 996 -660
rect 1360 -664 1756 -660
rect 2120 -664 2512 -660
rect 2516 -664 2520 -660
rect 2876 -664 3268 -660
rect 3272 -664 3276 -660
rect 240 -676 340 -672
rect 600 -984 996 -980
rect 1360 -984 1756 -980
rect 2120 -984 2512 -980
rect 2516 -984 2520 -980
rect 2876 -984 3268 -980
rect 3272 -984 3276 -980
rect 240 -992 340 -988
rect 1532 -1276 2228 -1272
rect 2320 -1276 3024 -1272
rect 44 -1280 748 -1276
rect 3056 -1284 3780 -1280
rect 768 -1288 1508 -1284
rect 2240 -1292 2432 -1288
rect 3028 -1292 3052 -1288
rect 2876 -1304 3268 -1300
rect 1278 -1352 1300 -1348
rect 2836 -1352 2852 -1348
rect 3784 -1364 3796 -1360
rect -88 -1484 -80 -1480
rect -76 -1484 -64 -1480
rect 2832 -1524 3796 -1520
rect 556 -1532 1300 -1528
rect 2028 -1544 2852 -1540
rect 1280 -1584 2016 -1580
<< m2contact >>
rect 236 288 240 292
rect 340 288 344 292
rect 748 288 752 292
rect 996 288 1000 292
rect 1508 288 1512 292
rect 1756 288 1760 292
rect 2268 288 2272 292
rect 2512 288 2516 292
rect 3024 288 3028 292
rect 3268 288 3272 292
rect 3780 288 3784 292
rect 596 -16 600 -12
rect 236 -32 240 -28
rect 340 -32 344 -28
rect 996 -16 1000 -12
rect 1356 -16 1360 -12
rect 1756 -16 1760 -12
rect 2116 -16 2120 -12
rect 2512 -16 2516 -12
rect 2872 -20 2876 -16
rect 3268 -20 3272 -16
rect 596 -340 600 -336
rect 236 -356 240 -352
rect 340 -356 344 -352
rect 996 -340 1000 -336
rect 1356 -340 1360 -336
rect 1756 -340 1760 -336
rect 2116 -340 2120 -336
rect 2512 -340 2516 -336
rect 2872 -340 2876 -336
rect 3268 -340 3272 -336
rect 596 -664 600 -660
rect 236 -676 240 -672
rect 340 -676 344 -672
rect 996 -664 1000 -660
rect 1356 -664 1360 -660
rect 1756 -664 1760 -660
rect 2116 -664 2120 -660
rect 2512 -664 2516 -660
rect 2872 -664 2876 -660
rect 3268 -664 3272 -660
rect 596 -984 600 -980
rect 236 -992 240 -988
rect 340 -992 344 -988
rect 996 -984 1000 -980
rect 1356 -984 1360 -980
rect 1756 -984 1760 -980
rect 2116 -984 2120 -980
rect 2512 -984 2516 -980
rect 2872 -984 2876 -980
rect 3268 -984 3272 -980
rect 364 -1224 368 -1220
rect 224 -1248 228 -1244
rect 40 -1280 44 -1276
rect 2684 -1224 2688 -1220
rect 596 -1260 600 -1256
rect 2228 -1264 2232 -1260
rect 748 -1280 752 -1276
rect 364 -1292 368 -1288
rect 764 -1288 768 -1284
rect 224 -1388 228 -1384
rect 552 -1420 556 -1416
rect -80 -1484 -76 -1480
rect 1508 -1288 1512 -1284
rect 1528 -1276 1532 -1272
rect 1100 -1304 1104 -1300
rect 916 -1400 920 -1396
rect 1300 -1352 1304 -1348
rect 552 -1532 556 -1528
rect 2228 -1276 2232 -1272
rect 2316 -1276 2320 -1272
rect 1860 -1292 1864 -1288
rect 1676 -1388 1680 -1384
rect 2016 -1340 2020 -1336
rect 1300 -1532 1304 -1528
rect 1276 -1584 1280 -1580
rect 2024 -1420 2028 -1416
rect 2236 -1292 2240 -1288
rect 2432 -1292 2436 -1288
rect 3648 -1224 3652 -1220
rect 3024 -1276 3028 -1272
rect 2684 -1304 2688 -1300
rect 3052 -1284 3056 -1280
rect 2872 -1304 2876 -1300
rect 3024 -1292 3028 -1288
rect 3052 -1292 3056 -1288
rect 2852 -1352 2856 -1348
rect 2828 -1432 2832 -1428
rect 2828 -1524 2832 -1520
rect 2024 -1544 2028 -1540
rect 3268 -1304 3272 -1300
rect 3780 -1284 3784 -1280
rect 3648 -1316 3652 -1312
rect 3796 -1364 3800 -1360
rect 3760 -1444 3764 -1440
rect 3796 -1524 3800 -1520
rect 2852 -1544 2856 -1540
rect 2016 -1584 2020 -1580
use adder2  adder2_1
timestamp 1607099119
transform 1 0 2208 0 1 -1464
box -28 -63 628 164
use multi  multi_4
timestamp 1607107347
transform 1 0 4 0 1 -1260
box -4 -40 3792 272
use adder2  adder2_0
timestamp 1607099119
transform 1 0 3160 0 1 -1476
box -28 -63 628 164
use adder2  adder2_2
timestamp 1607099119
transform 1 0 1404 0 1 -1452
box -28 -63 628 164
use adder2  adder2_3
timestamp 1607099119
transform 1 0 656 0 1 -1464
box -28 -63 628 164
use adder2  adder2_4
timestamp 1607099119
transform 1 0 -68 0 1 -1452
box -28 -63 628 164
use multi  multi_3
timestamp 1607107347
transform 1 0 4 0 1 -944
box -4 -40 3792 272
use multi  multi_2
timestamp 1607107347
transform 1 0 4 0 1 -624
box -4 -40 3792 272
use multi  multi_1
timestamp 1607107347
transform 1 0 4 0 1 -300
box -4 -40 3792 272
use multi  multi_0
timestamp 1607107347
transform 1 0 4 0 1 24
box -4 -40 3792 272
<< labels >>
rlabel metal1 3631 -18 3631 -18 1 p0
rlabel metal1 3631 -342 3631 -342 1 p1
rlabel metal1 3770 298 3770 298 5 a0
rlabel metal2 325 290 325 290 1 gnd
rlabel metal1 158 298 158 298 5 vdd
rlabel metal1 738 297 738 297 5 a4
rlabel metal1 1498 298 1498 298 5 a3
rlabel metal1 2258 298 2258 298 5 a2
rlabel metal1 3013 298 3013 298 5 a1
rlabel metal1 -2 94 -2 94 3 b0
rlabel metal1 -2 -230 -2 -230 3 b1
rlabel metal1 3631 -667 3631 -667 1 p2
rlabel metal1 3630 -986 3630 -986 1 p3
rlabel metal1 -2 -554 -2 -554 3 b2
rlabel metal1 -2 -874 -2 -874 3 b3
rlabel metal1 -1 -1190 -1 -1190 3 b4
rlabel metal1 3630 -1303 3630 -1303 1 p4
rlabel metal1 3482 -1538 3482 -1538 1 p5
rlabel metal1 2530 -1526 2530 -1526 1 p6
rlabel metal1 1726 -1514 1726 -1514 1 p7
rlabel metal1 978 -1526 978 -1526 1 p8
rlabel metal1 254 -1514 254 -1514 1 p9
<< end >>
