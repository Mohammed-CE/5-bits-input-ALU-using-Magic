magic
tech scmos
timestamp 1607190180
<< metal1 >>
rect 804 356 808 360
rect 428 220 432 224
rect 724 112 728 138
rect 1016 136 1020 140
rect 1016 108 1020 112
rect 1180 107 1184 141
rect 428 24 432 28
rect 752 -179 756 -24
rect 1308 -40 1312 288
rect 1320 248 1324 288
rect 1324 240 1328 244
rect 1336 4 1340 316
rect 1324 0 1340 4
rect 804 -112 808 -108
rect 892 -140 896 -120
rect 832 -156 836 -148
rect 1340 -216 1344 -44
rect 456 -288 460 -284
rect 752 -412 756 -345
rect 1044 -372 1048 -368
rect 1044 -400 1048 -396
rect 1208 -415 1212 -360
rect 456 -484 460 -480
rect 1332 -548 1336 -220
rect 1356 -264 1360 -72
rect 1372 -508 1376 -192
rect 1344 -512 1376 -508
rect 748 -661 752 -612
rect 832 -620 836 -616
rect 1204 -648 1208 -628
rect 828 -660 832 -656
rect 1332 -724 1336 -552
rect 1352 -768 1356 -580
rect 452 -796 456 -792
rect 1040 -880 1044 -876
<< metal2 >>
rect 1328 316 1336 320
rect 1320 -44 1340 -40
rect 1332 -72 1356 -68
rect 1356 -192 1372 -188
rect 1356 -700 1360 -696
<< m2contact >>
rect 1336 316 1340 320
rect 1308 288 1312 292
rect 752 -24 756 -20
rect 1320 288 1324 292
rect 1308 -44 1312 -40
rect 1340 -44 1344 -40
rect 892 -120 896 -116
rect 892 -144 896 -140
rect 1332 -220 1336 -216
rect 1340 -220 1344 -216
rect 1356 -72 1360 -68
rect 1372 -192 1376 -188
rect 1332 -552 1336 -548
rect 1204 -628 1208 -624
rect 1204 -652 1208 -648
rect 1332 -728 1336 -724
rect 1352 -580 1356 -576
use addsub  addsub_3
timestamp 1607190180
transform 1 0 680 0 -1 -416
box -220 -20 680 212
use addsub  addsub_0
timestamp 1607190180
transform 1 0 652 0 1 156
box -220 -20 680 212
use addsub  addsub_1
timestamp 1607190180
transform 1 0 652 0 -1 92
box -220 -20 680 212
use addsub  addsub_2
timestamp 1607190180
transform 1 0 680 0 1 -352
box -220 -20 680 212
use addsub  addsub_4
timestamp 1607190180
transform 1 0 676 0 1 -860
box -220 -20 680 212
<< end >>
