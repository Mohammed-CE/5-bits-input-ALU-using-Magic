magic
tech scmos
timestamp 1605560872
<< metal1 >>
rect 0 40 4 48
rect 0 -44 4 -36
<< metal2 >>
rect 0 96 4 100
rect 0 0 4 4
rect 0 -96 4 -92
<< m2contact >>
rect 0 48 4 52
rect 0 -48 4 -44
use not  not_1
timestamp 1605560378
transform 1 0 -36 0 -1 -48
box 4 -52 40 48
use not  not_0
timestamp 1605560378
transform 1 0 -36 0 1 52
box 4 -52 40 48
use and  and_1
timestamp 1605560441
transform 1 0 12 0 -1 4
box -12 0 68 100
use and  and_0
timestamp 1605560441
transform 1 0 12 0 1 0
box -12 0 68 100
<< end >>
